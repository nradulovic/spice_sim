* C:\Program Files (x86)\LTC\LTspiceIV\lib\sym\Draft1.asc
.subckt npn_therm 1 2 3 4
Q1 1 qb 3 0 {NPN}
B1 0 Pj I=IC(Q1)*V(1,3)
C1 Pj 0 {Cj}
R2 Pc Pj {Rjc}
C2 Pc 0 {Cc}
R3 4 Pc {Rch}
R4 4 0 90
E1 qb 2 Pj 0 {TCvbe}
.ends npn_therm
