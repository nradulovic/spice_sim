* Z:\home\nesa\Electronic\Active Projects\Simulation\Sims\LME49810.asc
Q1 5 N016 N022 0 NPN2
I1 3 N004 2.8m
Q2 3 N004 7 0 NPN2
Q3 4 5 8 0 PNP2
Q4 N004 N004 N005 0 NPN2
Q5 N005 N005 6 0 NPN2
C5 3 N004 6p
D1 5 6 zener
Q6 9 N015 N020 0 NPN1
Q7 N013 N015 N021 0 NPN1
R10 N021 4 10
R11 N020 4 10
Q8 9 N008 N006 0 PNP1
Q9 N013 N009 N007 0 PNP1
I2 3 N003 0.5m
C4 3 N003 5p
R13 3 N001 500k
R14 N003 N006 800
R15 N003 N007 800
V1 N009 N010 3m
Q10 3 2 N010 0 NPN1
Q11 3 1 N008 0 NPN1
Q12 N011 9 N016 0 NPN1
Q13 N011 N013 N015 0 NPN1
C10 N001 N003 1�
R9 N022 4 200
R16 3 N002 400k
C9 N002 N004 1�
Q14 vcc 0 N011 0 NPN1
Q15 N008 N014 N017 0 NPN1
Q16 N010 N014 N019 0 NPN1
R17 N019 4 39k
R18 N017 4 39k
Q17 N011 N012 N014 0 NPN1
R7 N011 N012 100k
V6 N018 4 2.5 Rser=1
D2 N012 N018 diode
Q18 N014 N024 N026 0 NPN1
Q19 N015 N024 N027 0 NPN1
Q20 N016 N024 N028 0 NPN1
R12 N027 4 5
R19 N028 4 5
R20 N026 4 5
Q21 N024 N024 N025 0 NPN1
R21 N025 4 5
I3 N011 N024 100�
R8 N011 N023 400k
C6 N023 N024 1�
.model npn1 npn (IS=2e-14 IKF=0.1 VAF=80 BF=320 RE=10 RB=50 RBM=1 IRB=50u CJC=3p CJE=8p XCJC=0.8)
.model npn2 npn (IS=2e-14 IKF=0.18 VAF=50 BF=150 RE=5 RB=100 RBM=7 IRB=20u CJC=6p CJE=9p XCJC=0.6)
.model pnp2 pnp (IS=2e-14 IKF=0.15 VAF=40 BF=100 RE=7 RB=150 RBM=10 IRB=20u CJC=7p CJE=10p XCJC=0.6)
.model pnp1 pnp (IS=2e-14 IKF=0.08 VAF=94 BF=250 RE=10 RB=70 RBM=2 IRB=50u CJC=4p CJE=9p)
.model diode D(Is=2.52n Rs=.568 N=1.752 Cjo=4p M=.4 tt=20n Iave=200m Vpk=75)
.model zener D(Is=.6n Rs=.5 Cjo=150p nbv=5 bv=10 Ibv=1m Vpk=10)
.end
